`timescale 1ns / 1ps
`default_nettype none
module  tone_detection_fsm(
            input wire clk_in,
            input wire rst_in,
            input wire [15:0] fft_data,
            output logic [3:0] tone_ident
  );
  
    

endmodule
`default_nettype wire

