`timescale 1ns / 1ps
`default_nettype none // prevents system from inferring an undeclared logic (good practice)
 
module top_level(
  input wire [15:0] sw, //all 16 input slide switches
  input wire [3:0] btn, //all four momentary button switches
  output logic [15:0] led, //16 green output LEDs (located right above switches)
  output logic [2:0] rgb0, //RGB channels of RGB LED0
  output logic [2:0] rgb1, //RGB channels of RGB LED1
  output logic [3:0] ss0_an,//anode control for upper four digits of seven-seg display
  output logic [3:0] ss1_an,//anode control for lower four digits of seven-seg display
  output logic [6:0] ss0_c, //cathode controls for the segments of upper four digits
  output logic [6:0] ss1_c //cathod controls for the segments of lower four digits
  );
 
  logic [6:0] ss0_cn, ss1_cn; //used for inverting output signal
 
  // instantiate a alu module called 'n1' that controls the upper four 7-seg
  alu n1(
    .d0_in(sw[7:0]),
    .d1_in(sw[15:8]),
    .sel_in(btn),
    .res_out(led[15:0]),
    .gt_out(rgb1[2]),
    .eq_out(rgb0[0])
      );

  assign {ss0_an, ss1_an} = 8'h01; // all low (on). to turn off digits, set high
  assign ss0_c = ~ss0_cn; //the cathodes on the seven segment are active low, so invert
  assign ss1_c = ~ss1_cn; //same as above
 
  /* we'll use the LEDs later...for now, just link them to the switches
   * and force some lights on
   */
 
  // assign led = sw;
  // assign rgb0[0] = 1'b1; //red channel of RGB LED 0
  // assign rgb1[2] = 1'b1; //blue channel of RGB LED 1

 
endmodule // top_level
/* I usually add a comment to associate my endmodule line with the module name
 * this helps when if you have multiple module definitions in a file
 */
 
// reset the default net type to wire, sometimes other code expects this.
`default_nettype wire